`define data_width 32
`define addr_width 32
`define no_of_transactions 200
